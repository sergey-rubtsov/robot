`define MODULE_NAME PWM_Top
`define WIDTH 10
